class agent_config extends uvm_object;
    `uvm_object_utils(agent_config)

    virtual conv_interface vif;
endclass